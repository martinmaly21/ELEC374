`timescale 1ns/ 1ps

module and_32_gate(
			input wire [31:0] a_in,
			input wire [31:0] b_in,
			output wire [31:0] c_out
			);
			
			
			genvar i;
			generate
					for(i = 0; i<32; i = i + 1)
						begin: gen_loop
							assign c_out[i] = ((a_in[i])&(b_in[i]));
						end
			endgenerate
endmodule
							
