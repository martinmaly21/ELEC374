

`timescale 1ns/10ps
module brmi_tb;

endmodule 