

`timescale 1ns/10ps
module brnz_tb;

endmodule 