

`timescale 1ns/10ps
module brpl_tb;

endmodule 