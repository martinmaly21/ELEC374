

`timescale 1ns/10ps
module brzr_tb;

endmodule 