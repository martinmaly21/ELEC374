module BUS ();

endmodule
